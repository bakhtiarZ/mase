module silu_lut(input logic [6:0] data_in_0, output logic [6:0] data_out_0);
    always_comb begin
        case(data_in_0)
            7'b0000000: data_out_0 = 7'b0000000;
            7'b0000001: data_out_0 = 7'b0000001;
            7'b0000010: data_out_0 = 7'b0000010;
            7'b0000011: data_out_0 = 7'b0000011;
            7'b0000100: data_out_0 = 7'b0000100;
            7'b0000101: data_out_0 = 7'b0000101;
            7'b0000110: data_out_0 = 7'b0000110;
            7'b0000111: data_out_0 = 7'b0000111;
            7'b0001000: data_out_0 = 7'b0001000;
            7'b0001001: data_out_0 = 7'b0001001;
            7'b0001010: data_out_0 = 7'b0001010;
            7'b0001011: data_out_0 = 7'b0001011;
            7'b0001100: data_out_0 = 7'b0001100;
            7'b0001101: data_out_0 = 7'b0001101;
            7'b0001110: data_out_0 = 7'b0001110;
            7'b0001111: data_out_0 = 7'b0001111;
            7'b0010000: data_out_0 = 7'b0010000;
            7'b0010001: data_out_0 = 7'b0010001;
            7'b0010010: data_out_0 = 7'b0010010;
            7'b0010011: data_out_0 = 7'b0010011;
            7'b0010100: data_out_0 = 7'b0010100;
            7'b0010101: data_out_0 = 7'b0010101;
            7'b0010110: data_out_0 = 7'b0010110;
            7'b0010111: data_out_0 = 7'b0010111;
            7'b0011000: data_out_0 = 7'b0011000;
            7'b0011001: data_out_0 = 7'b0011001;
            7'b0011010: data_out_0 = 7'b0011010;
            7'b0011011: data_out_0 = 7'b0011011;
            7'b0011100: data_out_0 = 7'b0011100;
            7'b0011101: data_out_0 = 7'b0011101;
            7'b0011110: data_out_0 = 7'b0011110;
            7'b0011111: data_out_0 = 7'b0011111;
            7'b0100000: data_out_0 = 7'b0100000;
            7'b0100001: data_out_0 = 7'b0100001;
            7'b0100010: data_out_0 = 7'b0100010;
            7'b0100011: data_out_0 = 7'b0100011;
            7'b0100100: data_out_0 = 7'b0100100;
            7'b0100101: data_out_0 = 7'b0100101;
            7'b0100110: data_out_0 = 7'b0100110;
            7'b0100111: data_out_0 = 7'b0100111;
            7'b0101000: data_out_0 = 7'b0101000;
            7'b0101001: data_out_0 = 7'b0101001;
            7'b0101010: data_out_0 = 7'b0101010;
            7'b0101011: data_out_0 = 7'b0101011;
            7'b0101100: data_out_0 = 7'b0101100;
            7'b0101101: data_out_0 = 7'b0101101;
            7'b0101110: data_out_0 = 7'b0101110;
            7'b0101111: data_out_0 = 7'b0101111;
            7'b0110000: data_out_0 = 7'b0110000;
            7'b0110001: data_out_0 = 7'b0110001;
            7'b0110010: data_out_0 = 7'b0110010;
            7'b0110011: data_out_0 = 7'b0110011;
            7'b0110100: data_out_0 = 7'b0110100;
            7'b0110101: data_out_0 = 7'b0110101;
            7'b0110110: data_out_0 = 7'b0110110;
            7'b0110111: data_out_0 = 7'b0110111;
            7'b0111000: data_out_0 = 7'b0111000;
            7'b0111001: data_out_0 = 7'b0111001;
            7'b0111010: data_out_0 = 7'b0111010;
            7'b0111011: data_out_0 = 7'b0111011;
            7'b0111100: data_out_0 = 7'b0111100;
            7'b0111101: data_out_0 = 7'b0111101;
            7'b0111110: data_out_0 = 7'b0111110;
            7'b0111111: data_out_0 = 7'b0111111;
            7'b1000000: data_out_0 = 7'b0000000;
            7'b1000001: data_out_0 = 7'b0000000;
            7'b1000010: data_out_0 = 7'b0000000;
            7'b1000011: data_out_0 = 7'b0000000;
            7'b1000100: data_out_0 = 7'b0000000;
            7'b1000101: data_out_0 = 7'b0000000;
            7'b1000110: data_out_0 = 7'b0000000;
            7'b1000111: data_out_0 = 7'b0000000;
            7'b1001000: data_out_0 = 7'b0000000;
            7'b1001001: data_out_0 = 7'b0000000;
            7'b1001010: data_out_0 = 7'b0000000;
            7'b1001011: data_out_0 = 7'b0000000;
            7'b1001100: data_out_0 = 7'b0000000;
            7'b1001101: data_out_0 = 7'b0000000;
            7'b1001110: data_out_0 = 7'b0000000;
            7'b1001111: data_out_0 = 7'b0000000;
            7'b1010000: data_out_0 = 7'b0000000;
            7'b1010001: data_out_0 = 7'b0000000;
            7'b1010010: data_out_0 = 7'b0000000;
            7'b1010011: data_out_0 = 7'b0000000;
            7'b1010100: data_out_0 = 7'b0000000;
            7'b1010101: data_out_0 = 7'b0000000;
            7'b1010110: data_out_0 = 7'b0000000;
            7'b1010111: data_out_0 = 7'b0000000;
            7'b1011000: data_out_0 = 7'b0000000;
            7'b1011001: data_out_0 = 7'b0000000;
            7'b1011010: data_out_0 = 7'b0000000;
            7'b1011011: data_out_0 = 7'b0000000;
            7'b1011100: data_out_0 = 7'b0000000;
            7'b1011101: data_out_0 = 7'b0000000;
            7'b1011110: data_out_0 = 7'b0000000;
            7'b1011111: data_out_0 = 7'b0000000;
            7'b1100000: data_out_0 = 7'b0000000;
            7'b1100001: data_out_0 = 7'b0000000;
            7'b1100010: data_out_0 = 7'b0000000;
            7'b1100011: data_out_0 = 7'b0000000;
            7'b1100100: data_out_0 = 7'b0000000;
            7'b1100101: data_out_0 = 7'b0000000;
            7'b1100110: data_out_0 = 7'b0000000;
            7'b1100111: data_out_0 = 7'b0000000;
            7'b1101000: data_out_0 = 7'b0000000;
            7'b1101001: data_out_0 = 7'b0000000;
            7'b1101010: data_out_0 = 7'b0000000;
            7'b1101011: data_out_0 = 7'b0000000;
            7'b1101100: data_out_0 = 7'b0000000;
            7'b1101101: data_out_0 = 7'b0000000;
            7'b1101110: data_out_0 = 7'b0000000;
            7'b1101111: data_out_0 = 7'b0000000;
            7'b1110000: data_out_0 = 7'b0000000;
            7'b1110001: data_out_0 = 7'b0000000;
            7'b1110010: data_out_0 = 7'b0000000;
            7'b1110011: data_out_0 = 7'b0000000;
            7'b1110100: data_out_0 = 7'b0000000;
            7'b1110101: data_out_0 = 7'b0000000;
            7'b1110110: data_out_0 = 7'b0000000;
            7'b1110111: data_out_0 = 7'b0000000;
            7'b1111000: data_out_0 = 7'b0000000;
            7'b1111001: data_out_0 = 7'b0000000;
            7'b1111010: data_out_0 = 7'b0000000;
            7'b1111011: data_out_0 = 7'b0000000;
            7'b1111100: data_out_0 = 7'b0000000;
            7'b1111101: data_out_0 = 7'b0000000;
            7'b1111110: data_out_0 = 7'b0000000;
            7'b1111111: data_out_0 = 7'b0000000;
            default: data_out_0 = 7'b0;
        endcase
    end
endmodule
