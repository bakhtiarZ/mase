module silu_lut(input logic [8:0] data_in_0, output logic [8:0] data_out_0);
    always_comb begin
        case(data_in_0)
            9'b000000000: data_out_0 = 9'b000000000;
            9'b000000001: data_out_0 = 9'b000000001;
            9'b000000010: data_out_0 = 9'b000000010;
            9'b000000011: data_out_0 = 9'b000000011;
            9'b000000100: data_out_0 = 9'b000000100;
            9'b000000101: data_out_0 = 9'b000000101;
            9'b000000110: data_out_0 = 9'b000000110;
            9'b000000111: data_out_0 = 9'b000000111;
            9'b000001000: data_out_0 = 9'b000001000;
            9'b000001001: data_out_0 = 9'b000001001;
            9'b000001010: data_out_0 = 9'b000001010;
            9'b000001011: data_out_0 = 9'b000001011;
            9'b000001100: data_out_0 = 9'b000001100;
            9'b000001101: data_out_0 = 9'b000001101;
            9'b000001110: data_out_0 = 9'b000001110;
            9'b000001111: data_out_0 = 9'b000001111;
            9'b000010000: data_out_0 = 9'b000010000;
            9'b000010001: data_out_0 = 9'b000010001;
            9'b000010010: data_out_0 = 9'b000010010;
            9'b000010011: data_out_0 = 9'b000010011;
            9'b000010100: data_out_0 = 9'b000010100;
            9'b000010101: data_out_0 = 9'b000010101;
            9'b000010110: data_out_0 = 9'b000010110;
            9'b000010111: data_out_0 = 9'b000010111;
            9'b000011000: data_out_0 = 9'b000011000;
            9'b000011001: data_out_0 = 9'b000011001;
            9'b000011010: data_out_0 = 9'b000011010;
            9'b000011011: data_out_0 = 9'b000011011;
            9'b000011100: data_out_0 = 9'b000011100;
            9'b000011101: data_out_0 = 9'b000011101;
            9'b000011110: data_out_0 = 9'b000011110;
            9'b000011111: data_out_0 = 9'b000011111;
            9'b000100000: data_out_0 = 9'b000100000;
            9'b000100001: data_out_0 = 9'b000100001;
            9'b000100010: data_out_0 = 9'b000100010;
            9'b000100011: data_out_0 = 9'b000100011;
            9'b000100100: data_out_0 = 9'b000100100;
            9'b000100101: data_out_0 = 9'b000100101;
            9'b000100110: data_out_0 = 9'b000100110;
            9'b000100111: data_out_0 = 9'b000100111;
            9'b000101000: data_out_0 = 9'b000101000;
            9'b000101001: data_out_0 = 9'b000101001;
            9'b000101010: data_out_0 = 9'b000101010;
            9'b000101011: data_out_0 = 9'b000101011;
            9'b000101100: data_out_0 = 9'b000101100;
            9'b000101101: data_out_0 = 9'b000101101;
            9'b000101110: data_out_0 = 9'b000101110;
            9'b000101111: data_out_0 = 9'b000101111;
            9'b000110000: data_out_0 = 9'b000110000;
            9'b000110001: data_out_0 = 9'b000110001;
            9'b000110010: data_out_0 = 9'b000110010;
            9'b000110011: data_out_0 = 9'b000110011;
            9'b000110100: data_out_0 = 9'b000110100;
            9'b000110101: data_out_0 = 9'b000110101;
            9'b000110110: data_out_0 = 9'b000110110;
            9'b000110111: data_out_0 = 9'b000110111;
            9'b000111000: data_out_0 = 9'b000111000;
            9'b000111001: data_out_0 = 9'b000111001;
            9'b000111010: data_out_0 = 9'b000111010;
            9'b000111011: data_out_0 = 9'b000111011;
            9'b000111100: data_out_0 = 9'b000111100;
            9'b000111101: data_out_0 = 9'b000111101;
            9'b000111110: data_out_0 = 9'b000111110;
            9'b000111111: data_out_0 = 9'b000111111;
            9'b001000000: data_out_0 = 9'b001000000;
            9'b001000001: data_out_0 = 9'b001000001;
            9'b001000010: data_out_0 = 9'b001000010;
            9'b001000011: data_out_0 = 9'b001000011;
            9'b001000100: data_out_0 = 9'b001000100;
            9'b001000101: data_out_0 = 9'b001000101;
            9'b001000110: data_out_0 = 9'b001000110;
            9'b001000111: data_out_0 = 9'b001000111;
            9'b001001000: data_out_0 = 9'b001001000;
            9'b001001001: data_out_0 = 9'b001001001;
            9'b001001010: data_out_0 = 9'b001001010;
            9'b001001011: data_out_0 = 9'b001001011;
            9'b001001100: data_out_0 = 9'b001001100;
            9'b001001101: data_out_0 = 9'b001001101;
            9'b001001110: data_out_0 = 9'b001001110;
            9'b001001111: data_out_0 = 9'b001001111;
            9'b001010000: data_out_0 = 9'b001010000;
            9'b001010001: data_out_0 = 9'b001010001;
            9'b001010010: data_out_0 = 9'b001010010;
            9'b001010011: data_out_0 = 9'b001010011;
            9'b001010100: data_out_0 = 9'b001010100;
            9'b001010101: data_out_0 = 9'b001010101;
            9'b001010110: data_out_0 = 9'b001010110;
            9'b001010111: data_out_0 = 9'b001010111;
            9'b001011000: data_out_0 = 9'b001011000;
            9'b001011001: data_out_0 = 9'b001011001;
            9'b001011010: data_out_0 = 9'b001011010;
            9'b001011011: data_out_0 = 9'b001011011;
            9'b001011100: data_out_0 = 9'b001011100;
            9'b001011101: data_out_0 = 9'b001011101;
            9'b001011110: data_out_0 = 9'b001011110;
            9'b001011111: data_out_0 = 9'b001011111;
            9'b001100000: data_out_0 = 9'b001100000;
            9'b001100001: data_out_0 = 9'b001100001;
            9'b001100010: data_out_0 = 9'b001100010;
            9'b001100011: data_out_0 = 9'b001100011;
            9'b001100100: data_out_0 = 9'b001100100;
            9'b001100101: data_out_0 = 9'b001100101;
            9'b001100110: data_out_0 = 9'b001100110;
            9'b001100111: data_out_0 = 9'b001100111;
            9'b001101000: data_out_0 = 9'b001101000;
            9'b001101001: data_out_0 = 9'b001101001;
            9'b001101010: data_out_0 = 9'b001101010;
            9'b001101011: data_out_0 = 9'b001101011;
            9'b001101100: data_out_0 = 9'b001101100;
            9'b001101101: data_out_0 = 9'b001101101;
            9'b001101110: data_out_0 = 9'b001101110;
            9'b001101111: data_out_0 = 9'b001101111;
            9'b001110000: data_out_0 = 9'b001110000;
            9'b001110001: data_out_0 = 9'b001110001;
            9'b001110010: data_out_0 = 9'b001110010;
            9'b001110011: data_out_0 = 9'b001110011;
            9'b001110100: data_out_0 = 9'b001110100;
            9'b001110101: data_out_0 = 9'b001110101;
            9'b001110110: data_out_0 = 9'b001110110;
            9'b001110111: data_out_0 = 9'b001110111;
            9'b001111000: data_out_0 = 9'b001111000;
            9'b001111001: data_out_0 = 9'b001111001;
            9'b001111010: data_out_0 = 9'b001111010;
            9'b001111011: data_out_0 = 9'b001111011;
            9'b001111100: data_out_0 = 9'b001111100;
            9'b001111101: data_out_0 = 9'b001111101;
            9'b001111110: data_out_0 = 9'b001111110;
            9'b001111111: data_out_0 = 9'b001111111;
            9'b010000000: data_out_0 = 9'b010000000;
            9'b010000001: data_out_0 = 9'b010000001;
            9'b010000010: data_out_0 = 9'b010000010;
            9'b010000011: data_out_0 = 9'b010000011;
            9'b010000100: data_out_0 = 9'b010000100;
            9'b010000101: data_out_0 = 9'b010000101;
            9'b010000110: data_out_0 = 9'b010000110;
            9'b010000111: data_out_0 = 9'b010000111;
            9'b010001000: data_out_0 = 9'b010001000;
            9'b010001001: data_out_0 = 9'b010001001;
            9'b010001010: data_out_0 = 9'b010001010;
            9'b010001011: data_out_0 = 9'b010001011;
            9'b010001100: data_out_0 = 9'b010001100;
            9'b010001101: data_out_0 = 9'b010001101;
            9'b010001110: data_out_0 = 9'b010001110;
            9'b010001111: data_out_0 = 9'b010001111;
            9'b010010000: data_out_0 = 9'b010010000;
            9'b010010001: data_out_0 = 9'b010010001;
            9'b010010010: data_out_0 = 9'b010010010;
            9'b010010011: data_out_0 = 9'b010010011;
            9'b010010100: data_out_0 = 9'b010010100;
            9'b010010101: data_out_0 = 9'b010010101;
            9'b010010110: data_out_0 = 9'b010010110;
            9'b010010111: data_out_0 = 9'b010010111;
            9'b010011000: data_out_0 = 9'b010011000;
            9'b010011001: data_out_0 = 9'b010011001;
            9'b010011010: data_out_0 = 9'b010011010;
            9'b010011011: data_out_0 = 9'b010011011;
            9'b010011100: data_out_0 = 9'b010011100;
            9'b010011101: data_out_0 = 9'b010011101;
            9'b010011110: data_out_0 = 9'b010011110;
            9'b010011111: data_out_0 = 9'b010011111;
            9'b010100000: data_out_0 = 9'b010100000;
            9'b010100001: data_out_0 = 9'b010100001;
            9'b010100010: data_out_0 = 9'b010100010;
            9'b010100011: data_out_0 = 9'b010100011;
            9'b010100100: data_out_0 = 9'b010100100;
            9'b010100101: data_out_0 = 9'b010100101;
            9'b010100110: data_out_0 = 9'b010100110;
            9'b010100111: data_out_0 = 9'b010100111;
            9'b010101000: data_out_0 = 9'b010101000;
            9'b010101001: data_out_0 = 9'b010101001;
            9'b010101010: data_out_0 = 9'b010101010;
            9'b010101011: data_out_0 = 9'b010101011;
            9'b010101100: data_out_0 = 9'b010101100;
            9'b010101101: data_out_0 = 9'b010101101;
            9'b010101110: data_out_0 = 9'b010101110;
            9'b010101111: data_out_0 = 9'b010101111;
            9'b010110000: data_out_0 = 9'b010110000;
            9'b010110001: data_out_0 = 9'b010110001;
            9'b010110010: data_out_0 = 9'b010110010;
            9'b010110011: data_out_0 = 9'b010110011;
            9'b010110100: data_out_0 = 9'b010110100;
            9'b010110101: data_out_0 = 9'b010110101;
            9'b010110110: data_out_0 = 9'b010110110;
            9'b010110111: data_out_0 = 9'b010110111;
            9'b010111000: data_out_0 = 9'b010111000;
            9'b010111001: data_out_0 = 9'b010111001;
            9'b010111010: data_out_0 = 9'b010111010;
            9'b010111011: data_out_0 = 9'b010111011;
            9'b010111100: data_out_0 = 9'b010111100;
            9'b010111101: data_out_0 = 9'b010111101;
            9'b010111110: data_out_0 = 9'b010111110;
            9'b010111111: data_out_0 = 9'b010111111;
            9'b011000000: data_out_0 = 9'b011000000;
            9'b011000001: data_out_0 = 9'b011000001;
            9'b011000010: data_out_0 = 9'b011000010;
            9'b011000011: data_out_0 = 9'b011000011;
            9'b011000100: data_out_0 = 9'b011000100;
            9'b011000101: data_out_0 = 9'b011000101;
            9'b011000110: data_out_0 = 9'b011000110;
            9'b011000111: data_out_0 = 9'b011000111;
            9'b011001000: data_out_0 = 9'b011001000;
            9'b011001001: data_out_0 = 9'b011001001;
            9'b011001010: data_out_0 = 9'b011001010;
            9'b011001011: data_out_0 = 9'b011001011;
            9'b011001100: data_out_0 = 9'b011001100;
            9'b011001101: data_out_0 = 9'b011001101;
            9'b011001110: data_out_0 = 9'b011001110;
            9'b011001111: data_out_0 = 9'b011001111;
            9'b011010000: data_out_0 = 9'b011010000;
            9'b011010001: data_out_0 = 9'b011010001;
            9'b011010010: data_out_0 = 9'b011010010;
            9'b011010011: data_out_0 = 9'b011010011;
            9'b011010100: data_out_0 = 9'b011010100;
            9'b011010101: data_out_0 = 9'b011010101;
            9'b011010110: data_out_0 = 9'b011010110;
            9'b011010111: data_out_0 = 9'b011010111;
            9'b011011000: data_out_0 = 9'b011011000;
            9'b011011001: data_out_0 = 9'b011011001;
            9'b011011010: data_out_0 = 9'b011011010;
            9'b011011011: data_out_0 = 9'b011011011;
            9'b011011100: data_out_0 = 9'b011011100;
            9'b011011101: data_out_0 = 9'b011011101;
            9'b011011110: data_out_0 = 9'b011011110;
            9'b011011111: data_out_0 = 9'b011011111;
            9'b011100000: data_out_0 = 9'b011100000;
            9'b011100001: data_out_0 = 9'b011100001;
            9'b011100010: data_out_0 = 9'b011100010;
            9'b011100011: data_out_0 = 9'b011100011;
            9'b011100100: data_out_0 = 9'b011100100;
            9'b011100101: data_out_0 = 9'b011100101;
            9'b011100110: data_out_0 = 9'b011100110;
            9'b011100111: data_out_0 = 9'b011100111;
            9'b011101000: data_out_0 = 9'b011101000;
            9'b011101001: data_out_0 = 9'b011101001;
            9'b011101010: data_out_0 = 9'b011101010;
            9'b011101011: data_out_0 = 9'b011101011;
            9'b011101100: data_out_0 = 9'b011101100;
            9'b011101101: data_out_0 = 9'b011101101;
            9'b011101110: data_out_0 = 9'b011101110;
            9'b011101111: data_out_0 = 9'b011101111;
            9'b011110000: data_out_0 = 9'b011110000;
            9'b011110001: data_out_0 = 9'b011110001;
            9'b011110010: data_out_0 = 9'b011110010;
            9'b011110011: data_out_0 = 9'b011110011;
            9'b011110100: data_out_0 = 9'b011110100;
            9'b011110101: data_out_0 = 9'b011110101;
            9'b011110110: data_out_0 = 9'b011110110;
            9'b011110111: data_out_0 = 9'b011110111;
            9'b011111000: data_out_0 = 9'b011111000;
            9'b011111001: data_out_0 = 9'b011111001;
            9'b011111010: data_out_0 = 9'b011111010;
            9'b011111011: data_out_0 = 9'b011111011;
            9'b011111100: data_out_0 = 9'b011111100;
            9'b011111101: data_out_0 = 9'b011111101;
            9'b011111110: data_out_0 = 9'b011111110;
            9'b011111111: data_out_0 = 9'b011111111;
            9'b100000000: data_out_0 = 9'b000000000;
            9'b100000001: data_out_0 = 9'b000000000;
            9'b100000010: data_out_0 = 9'b000000000;
            9'b100000011: data_out_0 = 9'b000000000;
            9'b100000100: data_out_0 = 9'b000000000;
            9'b100000101: data_out_0 = 9'b000000000;
            9'b100000110: data_out_0 = 9'b000000000;
            9'b100000111: data_out_0 = 9'b000000000;
            9'b100001000: data_out_0 = 9'b000000000;
            9'b100001001: data_out_0 = 9'b000000000;
            9'b100001010: data_out_0 = 9'b000000000;
            9'b100001011: data_out_0 = 9'b000000000;
            9'b100001100: data_out_0 = 9'b000000000;
            9'b100001101: data_out_0 = 9'b000000000;
            9'b100001110: data_out_0 = 9'b000000000;
            9'b100001111: data_out_0 = 9'b000000000;
            9'b100010000: data_out_0 = 9'b000000000;
            9'b100010001: data_out_0 = 9'b000000000;
            9'b100010010: data_out_0 = 9'b000000000;
            9'b100010011: data_out_0 = 9'b000000000;
            9'b100010100: data_out_0 = 9'b000000000;
            9'b100010101: data_out_0 = 9'b000000000;
            9'b100010110: data_out_0 = 9'b000000000;
            9'b100010111: data_out_0 = 9'b000000000;
            9'b100011000: data_out_0 = 9'b000000000;
            9'b100011001: data_out_0 = 9'b000000000;
            9'b100011010: data_out_0 = 9'b000000000;
            9'b100011011: data_out_0 = 9'b000000000;
            9'b100011100: data_out_0 = 9'b000000000;
            9'b100011101: data_out_0 = 9'b000000000;
            9'b100011110: data_out_0 = 9'b000000000;
            9'b100011111: data_out_0 = 9'b000000000;
            9'b100100000: data_out_0 = 9'b000000000;
            9'b100100001: data_out_0 = 9'b000000000;
            9'b100100010: data_out_0 = 9'b000000000;
            9'b100100011: data_out_0 = 9'b000000000;
            9'b100100100: data_out_0 = 9'b000000000;
            9'b100100101: data_out_0 = 9'b000000000;
            9'b100100110: data_out_0 = 9'b000000000;
            9'b100100111: data_out_0 = 9'b000000000;
            9'b100101000: data_out_0 = 9'b000000000;
            9'b100101001: data_out_0 = 9'b000000000;
            9'b100101010: data_out_0 = 9'b000000000;
            9'b100101011: data_out_0 = 9'b000000000;
            9'b100101100: data_out_0 = 9'b000000000;
            9'b100101101: data_out_0 = 9'b000000000;
            9'b100101110: data_out_0 = 9'b000000000;
            9'b100101111: data_out_0 = 9'b000000000;
            9'b100110000: data_out_0 = 9'b000000000;
            9'b100110001: data_out_0 = 9'b000000000;
            9'b100110010: data_out_0 = 9'b000000000;
            9'b100110011: data_out_0 = 9'b000000000;
            9'b100110100: data_out_0 = 9'b000000000;
            9'b100110101: data_out_0 = 9'b000000000;
            9'b100110110: data_out_0 = 9'b000000000;
            9'b100110111: data_out_0 = 9'b000000000;
            9'b100111000: data_out_0 = 9'b000000000;
            9'b100111001: data_out_0 = 9'b000000000;
            9'b100111010: data_out_0 = 9'b000000000;
            9'b100111011: data_out_0 = 9'b000000000;
            9'b100111100: data_out_0 = 9'b000000000;
            9'b100111101: data_out_0 = 9'b000000000;
            9'b100111110: data_out_0 = 9'b000000000;
            9'b100111111: data_out_0 = 9'b000000000;
            9'b101000000: data_out_0 = 9'b000000000;
            9'b101000001: data_out_0 = 9'b000000000;
            9'b101000010: data_out_0 = 9'b000000000;
            9'b101000011: data_out_0 = 9'b000000000;
            9'b101000100: data_out_0 = 9'b000000000;
            9'b101000101: data_out_0 = 9'b000000000;
            9'b101000110: data_out_0 = 9'b000000000;
            9'b101000111: data_out_0 = 9'b000000000;
            9'b101001000: data_out_0 = 9'b000000000;
            9'b101001001: data_out_0 = 9'b000000000;
            9'b101001010: data_out_0 = 9'b000000000;
            9'b101001011: data_out_0 = 9'b000000000;
            9'b101001100: data_out_0 = 9'b000000000;
            9'b101001101: data_out_0 = 9'b000000000;
            9'b101001110: data_out_0 = 9'b000000000;
            9'b101001111: data_out_0 = 9'b000000000;
            9'b101010000: data_out_0 = 9'b000000000;
            9'b101010001: data_out_0 = 9'b000000000;
            9'b101010010: data_out_0 = 9'b000000000;
            9'b101010011: data_out_0 = 9'b000000000;
            9'b101010100: data_out_0 = 9'b000000000;
            9'b101010101: data_out_0 = 9'b000000000;
            9'b101010110: data_out_0 = 9'b000000000;
            9'b101010111: data_out_0 = 9'b000000000;
            9'b101011000: data_out_0 = 9'b000000000;
            9'b101011001: data_out_0 = 9'b000000000;
            9'b101011010: data_out_0 = 9'b000000000;
            9'b101011011: data_out_0 = 9'b000000000;
            9'b101011100: data_out_0 = 9'b000000000;
            9'b101011101: data_out_0 = 9'b000000000;
            9'b101011110: data_out_0 = 9'b000000000;
            9'b101011111: data_out_0 = 9'b000000000;
            9'b101100000: data_out_0 = 9'b000000000;
            9'b101100001: data_out_0 = 9'b000000000;
            9'b101100010: data_out_0 = 9'b000000000;
            9'b101100011: data_out_0 = 9'b000000000;
            9'b101100100: data_out_0 = 9'b000000000;
            9'b101100101: data_out_0 = 9'b000000000;
            9'b101100110: data_out_0 = 9'b000000000;
            9'b101100111: data_out_0 = 9'b000000000;
            9'b101101000: data_out_0 = 9'b000000000;
            9'b101101001: data_out_0 = 9'b000000000;
            9'b101101010: data_out_0 = 9'b000000000;
            9'b101101011: data_out_0 = 9'b000000000;
            9'b101101100: data_out_0 = 9'b000000000;
            9'b101101101: data_out_0 = 9'b000000000;
            9'b101101110: data_out_0 = 9'b000000000;
            9'b101101111: data_out_0 = 9'b000000000;
            9'b101110000: data_out_0 = 9'b000000000;
            9'b101110001: data_out_0 = 9'b000000000;
            9'b101110010: data_out_0 = 9'b000000000;
            9'b101110011: data_out_0 = 9'b000000000;
            9'b101110100: data_out_0 = 9'b000000000;
            9'b101110101: data_out_0 = 9'b000000000;
            9'b101110110: data_out_0 = 9'b000000000;
            9'b101110111: data_out_0 = 9'b000000000;
            9'b101111000: data_out_0 = 9'b000000000;
            9'b101111001: data_out_0 = 9'b000000000;
            9'b101111010: data_out_0 = 9'b000000000;
            9'b101111011: data_out_0 = 9'b000000000;
            9'b101111100: data_out_0 = 9'b000000000;
            9'b101111101: data_out_0 = 9'b000000000;
            9'b101111110: data_out_0 = 9'b000000000;
            9'b101111111: data_out_0 = 9'b000000000;
            9'b110000000: data_out_0 = 9'b000000000;
            9'b110000001: data_out_0 = 9'b000000000;
            9'b110000010: data_out_0 = 9'b000000000;
            9'b110000011: data_out_0 = 9'b000000000;
            9'b110000100: data_out_0 = 9'b000000000;
            9'b110000101: data_out_0 = 9'b000000000;
            9'b110000110: data_out_0 = 9'b000000000;
            9'b110000111: data_out_0 = 9'b000000000;
            9'b110001000: data_out_0 = 9'b000000000;
            9'b110001001: data_out_0 = 9'b000000000;
            9'b110001010: data_out_0 = 9'b000000000;
            9'b110001011: data_out_0 = 9'b000000000;
            9'b110001100: data_out_0 = 9'b000000000;
            9'b110001101: data_out_0 = 9'b000000000;
            9'b110001110: data_out_0 = 9'b000000000;
            9'b110001111: data_out_0 = 9'b000000000;
            9'b110010000: data_out_0 = 9'b000000000;
            9'b110010001: data_out_0 = 9'b000000000;
            9'b110010010: data_out_0 = 9'b000000000;
            9'b110010011: data_out_0 = 9'b000000000;
            9'b110010100: data_out_0 = 9'b000000000;
            9'b110010101: data_out_0 = 9'b000000000;
            9'b110010110: data_out_0 = 9'b000000000;
            9'b110010111: data_out_0 = 9'b000000000;
            9'b110011000: data_out_0 = 9'b000000000;
            9'b110011001: data_out_0 = 9'b000000000;
            9'b110011010: data_out_0 = 9'b000000000;
            9'b110011011: data_out_0 = 9'b000000000;
            9'b110011100: data_out_0 = 9'b000000000;
            9'b110011101: data_out_0 = 9'b000000000;
            9'b110011110: data_out_0 = 9'b000000000;
            9'b110011111: data_out_0 = 9'b000000000;
            9'b110100000: data_out_0 = 9'b000000000;
            9'b110100001: data_out_0 = 9'b000000000;
            9'b110100010: data_out_0 = 9'b000000000;
            9'b110100011: data_out_0 = 9'b000000000;
            9'b110100100: data_out_0 = 9'b000000000;
            9'b110100101: data_out_0 = 9'b000000000;
            9'b110100110: data_out_0 = 9'b000000000;
            9'b110100111: data_out_0 = 9'b000000000;
            9'b110101000: data_out_0 = 9'b000000000;
            9'b110101001: data_out_0 = 9'b000000000;
            9'b110101010: data_out_0 = 9'b000000000;
            9'b110101011: data_out_0 = 9'b000000000;
            9'b110101100: data_out_0 = 9'b000000000;
            9'b110101101: data_out_0 = 9'b000000000;
            9'b110101110: data_out_0 = 9'b000000000;
            9'b110101111: data_out_0 = 9'b000000000;
            9'b110110000: data_out_0 = 9'b000000000;
            9'b110110001: data_out_0 = 9'b000000000;
            9'b110110010: data_out_0 = 9'b000000000;
            9'b110110011: data_out_0 = 9'b000000000;
            9'b110110100: data_out_0 = 9'b000000000;
            9'b110110101: data_out_0 = 9'b000000000;
            9'b110110110: data_out_0 = 9'b000000000;
            9'b110110111: data_out_0 = 9'b000000000;
            9'b110111000: data_out_0 = 9'b000000000;
            9'b110111001: data_out_0 = 9'b000000000;
            9'b110111010: data_out_0 = 9'b000000000;
            9'b110111011: data_out_0 = 9'b000000000;
            9'b110111100: data_out_0 = 9'b000000000;
            9'b110111101: data_out_0 = 9'b000000000;
            9'b110111110: data_out_0 = 9'b000000000;
            9'b110111111: data_out_0 = 9'b000000000;
            9'b111000000: data_out_0 = 9'b000000000;
            9'b111000001: data_out_0 = 9'b000000000;
            9'b111000010: data_out_0 = 9'b000000000;
            9'b111000011: data_out_0 = 9'b000000000;
            9'b111000100: data_out_0 = 9'b000000000;
            9'b111000101: data_out_0 = 9'b000000000;
            9'b111000110: data_out_0 = 9'b000000000;
            9'b111000111: data_out_0 = 9'b000000000;
            9'b111001000: data_out_0 = 9'b000000000;
            9'b111001001: data_out_0 = 9'b000000000;
            9'b111001010: data_out_0 = 9'b000000000;
            9'b111001011: data_out_0 = 9'b000000000;
            9'b111001100: data_out_0 = 9'b000000000;
            9'b111001101: data_out_0 = 9'b000000000;
            9'b111001110: data_out_0 = 9'b000000000;
            9'b111001111: data_out_0 = 9'b000000000;
            9'b111010000: data_out_0 = 9'b000000000;
            9'b111010001: data_out_0 = 9'b000000000;
            9'b111010010: data_out_0 = 9'b000000000;
            9'b111010011: data_out_0 = 9'b000000000;
            9'b111010100: data_out_0 = 9'b000000000;
            9'b111010101: data_out_0 = 9'b000000000;
            9'b111010110: data_out_0 = 9'b000000000;
            9'b111010111: data_out_0 = 9'b000000000;
            9'b111011000: data_out_0 = 9'b000000000;
            9'b111011001: data_out_0 = 9'b000000000;
            9'b111011010: data_out_0 = 9'b000000000;
            9'b111011011: data_out_0 = 9'b000000000;
            9'b111011100: data_out_0 = 9'b000000000;
            9'b111011101: data_out_0 = 9'b000000000;
            9'b111011110: data_out_0 = 9'b000000000;
            9'b111011111: data_out_0 = 9'b000000000;
            9'b111100000: data_out_0 = 9'b000000000;
            9'b111100001: data_out_0 = 9'b000000000;
            9'b111100010: data_out_0 = 9'b000000000;
            9'b111100011: data_out_0 = 9'b000000000;
            9'b111100100: data_out_0 = 9'b000000000;
            9'b111100101: data_out_0 = 9'b000000000;
            9'b111100110: data_out_0 = 9'b000000000;
            9'b111100111: data_out_0 = 9'b000000000;
            9'b111101000: data_out_0 = 9'b000000000;
            9'b111101001: data_out_0 = 9'b000000000;
            9'b111101010: data_out_0 = 9'b000000000;
            9'b111101011: data_out_0 = 9'b000000000;
            9'b111101100: data_out_0 = 9'b000000000;
            9'b111101101: data_out_0 = 9'b000000000;
            9'b111101110: data_out_0 = 9'b000000000;
            9'b111101111: data_out_0 = 9'b000000000;
            9'b111110000: data_out_0 = 9'b000000000;
            9'b111110001: data_out_0 = 9'b000000000;
            9'b111110010: data_out_0 = 9'b000000000;
            9'b111110011: data_out_0 = 9'b000000000;
            9'b111110100: data_out_0 = 9'b000000000;
            9'b111110101: data_out_0 = 9'b000000000;
            9'b111110110: data_out_0 = 9'b000000000;
            9'b111110111: data_out_0 = 9'b000000000;
            9'b111111000: data_out_0 = 9'b000000000;
            9'b111111001: data_out_0 = 9'b000000000;
            9'b111111010: data_out_0 = 9'b000000000;
            9'b111111011: data_out_0 = 9'b000000000;
            9'b111111100: data_out_0 = 9'b000000000;
            9'b111111101: data_out_0 = 9'b000000000;
            9'b111111110: data_out_0 = 9'b000000000;
            9'b111111111: data_out_0 = 9'b000000000;
            default: data_out_0 = 9'b0;
        endcase
    end
endmodule
